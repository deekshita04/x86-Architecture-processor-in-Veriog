

module and_vector(output [63:0] Y, input [63:0] A ,input [63:0] B, output overflow);

  assign overflow = 0;
  genvar i;
  generate
    for(i=0 ; i<64 ; i=i+1)
    begin
      and gate(Y[i],A[i],B[i]);
    end
  endgenerate
endmodule

//`timescale 1ns / 1ps
//module tb_AND_block_64;
//  reg [63:0] A, B;
//  wire [63:0] Y;
//  AND_block_64 uut (
//    .Y(Y),
//    .A(A),
//    .B(B)
//  );
//  initial begin
//    $dumpfile("and_block.vcd");
//    $dumpvars(0, tb_AND_block_64);
//        A = 64'b1101101101101101101101101101101101101101101101101101101101101101;
//        B = 64'b0010101010101010101010101010101010101010101010101010101010101010;
//        $monitor("Test Case 1: A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        A = 64'b1101101101101101101101101101101101101101101101101101101101101101;
//        B = 64'b1010101010101010101010101010101010101010101010101010101010101010;
//        $monitor("Test Case 2:A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        A = 64'b0111001110011100111001110011100111001110011100111001110011100;
//        B = 64'b1000111100001111000011110000111100001111000011110000111100000;
//        $monitor("Test Case 3:A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        A = 64'b0111001110011100111001110011100111001110011100111001110011100;
//        B = 64'b1000111100001111000011110000111100001111000011110000111100000;
//        $monitor("Test Case 4: A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        A = 64'b1111111111111111111111111111111111111111111111111111111111111110;
//        B = 64'b1111111111111111111111111111111111111111111111111111111111111110;
//        $monitor("Test Case 5: A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        A = 64'b0111111111111111111111111111111111111111111111111111111111111111;
//        B = 64'b0111111111111111111111111111111111111111111111111111111111111111;
//        $monitor("Test Case 6: A=%b, B=%b,Y=%b",A,B,Y);
//        #10
//        $finish;
//  end
//
//endmodule
//
//
//
//